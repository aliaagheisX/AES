module Shift_Rows_tb;
reg [127:0]in;
reg clk;
wire [127:0]out;

initial begin
clk = 0;
in = 128'hd42711aee0bf98f1b8b45de51e415230;
end

always #40 clk=~clk;


Shift_Rows uut(.in(in),.out(out),.clk(clk));
endmodule

/* 
d4e0b81e27bfb44111985d52aef1e530*/